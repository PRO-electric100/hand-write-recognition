library verilog;
use verilog.vl_types.all;
entity ALU_EXT_vlg_vec_tst is
end ALU_EXT_vlg_vec_tst;
